library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity NOR_Gate is
    Port (
        A : in STD_LOGIC;
        B : in STD_LOGIC;
        Y : out STD_LOGIC
    );
end NOR_Gate;

architecture Behavioral of NOR_Gate is
begin
    Y <= not (A or B);
end Behavioral;
